module ();

  initial
    begin

    end
  
endmodule

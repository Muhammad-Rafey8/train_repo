module ();
LOGIC a;
Logic b;
  initial
    begin

    end
  
endmodule

module ();
LOGIC a;
  initial
    begin

    end
  
endmodule
